-- Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, the Altera Quartus II License Agreement,
-- the Altera MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Altera and sold by Altera or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 15.0.1 Build 150 06/03/2015 SJ Web Edition"
-- CREATED		"Sun Oct 11 21:58:42 2015"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY sub3 IS 
	PORT
	(
		delayIN :  IN  STD_LOGIC;
		delayEN :  IN  STD_LOGIC;
		n3 :  OUT  STD_LOGIC;
		n4 :  OUT  STD_LOGIC;
		n5 :  OUT  STD_LOGIC;
		n6 :  OUT  STD_LOGIC;
		n7 :  OUT  STD_LOGIC;
		n8 :  OUT  STD_LOGIC;
		n9 :  OUT  STD_LOGIC;
		n10 :  OUT  STD_LOGIC;
		n11 :  OUT  STD_LOGIC;
		n12 :  OUT  STD_LOGIC;
		n13 :  OUT  STD_LOGIC;
		n14 :  OUT  STD_LOGIC;
		n15 :  OUT  STD_LOGIC;
		n16 :  OUT  STD_LOGIC;
		n17 :  OUT  STD_LOGIC;
		n18 :  OUT  STD_LOGIC;
		n19 :  OUT  STD_LOGIC;
		n20 :  OUT  STD_LOGIC;
		n21 :  OUT  STD_LOGIC;
		n22 :  OUT  STD_LOGIC;
		ENOout :  OUT  STD_LOGIC;
		INOout :  OUT  STD_LOGIC
	);
END sub3;

ARCHITECTURE bdf_type OF sub3 IS 

COMPONENT delaycellv3
	PORT(ENp : IN STD_LOGIC;
		 Reset : IN STD_LOGIC;
		 dIN : IN STD_LOGIC;
		 ENOp : OUT STD_LOGIC;
		 dOUT : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;


BEGIN 
n3 <= SYNTHESIZED_WIRE_2;
n4 <= SYNTHESIZED_WIRE_60;
n5 <= SYNTHESIZED_WIRE_58;
n6 <= SYNTHESIZED_WIRE_59;
n7 <= SYNTHESIZED_WIRE_61;
n8 <= SYNTHESIZED_WIRE_62;
n9 <= SYNTHESIZED_WIRE_63;
n10 <= SYNTHESIZED_WIRE_64;
n11 <= SYNTHESIZED_WIRE_65;
n12 <= SYNTHESIZED_WIRE_66;
n13 <= SYNTHESIZED_WIRE_67;
n14 <= SYNTHESIZED_WIRE_68;
n15 <= SYNTHESIZED_WIRE_69;
n16 <= SYNTHESIZED_WIRE_70;
n17 <= SYNTHESIZED_WIRE_71;
n18 <= SYNTHESIZED_WIRE_72;
n19 <= SYNTHESIZED_WIRE_73;
n20 <= SYNTHESIZED_WIRE_74;
n21 <= SYNTHESIZED_WIRE_75;
n22 <= SYNTHESIZED_WIRE_76;
INOout <= SYNTHESIZED_WIRE_76;



b2v_inst19 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_0,
		 Reset => SYNTHESIZED_WIRE_58,
		 dIN => SYNTHESIZED_WIRE_2,
		 ENOp => SYNTHESIZED_WIRE_3,
		 dOUT => SYNTHESIZED_WIRE_60);


b2v_inst23 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_3,
		 Reset => SYNTHESIZED_WIRE_59,
		 dIN => SYNTHESIZED_WIRE_60,
		 ENOp => SYNTHESIZED_WIRE_6,
		 dOUT => SYNTHESIZED_WIRE_58);


b2v_inst24 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_6,
		 Reset => SYNTHESIZED_WIRE_61,
		 dIN => SYNTHESIZED_WIRE_58,
		 ENOp => SYNTHESIZED_WIRE_9,
		 dOUT => SYNTHESIZED_WIRE_59);


b2v_inst25 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_9,
		 Reset => SYNTHESIZED_WIRE_62,
		 dIN => SYNTHESIZED_WIRE_59,
		 ENOp => SYNTHESIZED_WIRE_12,
		 dOUT => SYNTHESIZED_WIRE_61);


b2v_inst26 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_12,
		 Reset => SYNTHESIZED_WIRE_63,
		 dIN => SYNTHESIZED_WIRE_61,
		 ENOp => SYNTHESIZED_WIRE_15,
		 dOUT => SYNTHESIZED_WIRE_62);


b2v_inst27 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_15,
		 Reset => SYNTHESIZED_WIRE_64,
		 dIN => SYNTHESIZED_WIRE_62,
		 ENOp => SYNTHESIZED_WIRE_19,
		 dOUT => SYNTHESIZED_WIRE_63);


b2v_inst28 : delaycellv3
PORT MAP(ENp => delayEN,
		 Reset => SYNTHESIZED_WIRE_60,
		 dIN => delayIN,
		 ENOp => SYNTHESIZED_WIRE_0,
		 dOUT => SYNTHESIZED_WIRE_2);


b2v_inst29 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_19,
		 Reset => SYNTHESIZED_WIRE_65,
		 dIN => SYNTHESIZED_WIRE_63,
		 ENOp => SYNTHESIZED_WIRE_22,
		 dOUT => SYNTHESIZED_WIRE_64);


b2v_inst30 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_22,
		 Reset => SYNTHESIZED_WIRE_66,
		 dIN => SYNTHESIZED_WIRE_64,
		 ENOp => SYNTHESIZED_WIRE_25,
		 dOUT => SYNTHESIZED_WIRE_65);


b2v_inst31 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_25,
		 Reset => SYNTHESIZED_WIRE_67,
		 dIN => SYNTHESIZED_WIRE_65,
		 ENOp => SYNTHESIZED_WIRE_28,
		 dOUT => SYNTHESIZED_WIRE_66);


b2v_inst32 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_28,
		 Reset => SYNTHESIZED_WIRE_68,
		 dIN => SYNTHESIZED_WIRE_66,
		 ENOp => SYNTHESIZED_WIRE_31,
		 dOUT => SYNTHESIZED_WIRE_67);


b2v_inst33 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_31,
		 Reset => SYNTHESIZED_WIRE_69,
		 dIN => SYNTHESIZED_WIRE_67,
		 ENOp => SYNTHESIZED_WIRE_34,
		 dOUT => SYNTHESIZED_WIRE_68);


b2v_inst34 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_34,
		 Reset => SYNTHESIZED_WIRE_70,
		 dIN => SYNTHESIZED_WIRE_68,
		 ENOp => SYNTHESIZED_WIRE_37,
		 dOUT => SYNTHESIZED_WIRE_69);


b2v_inst35 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_37,
		 Reset => SYNTHESIZED_WIRE_71,
		 dIN => SYNTHESIZED_WIRE_69,
		 ENOp => SYNTHESIZED_WIRE_40,
		 dOUT => SYNTHESIZED_WIRE_70);


b2v_inst36 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_40,
		 Reset => SYNTHESIZED_WIRE_72,
		 dIN => SYNTHESIZED_WIRE_70,
		 ENOp => SYNTHESIZED_WIRE_43,
		 dOUT => SYNTHESIZED_WIRE_71);


b2v_inst37 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_43,
		 Reset => SYNTHESIZED_WIRE_73,
		 dIN => SYNTHESIZED_WIRE_71,
		 ENOp => SYNTHESIZED_WIRE_46,
		 dOUT => SYNTHESIZED_WIRE_72);


b2v_inst38 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_46,
		 Reset => SYNTHESIZED_WIRE_74,
		 dIN => SYNTHESIZED_WIRE_72,
		 ENOp => SYNTHESIZED_WIRE_49,
		 dOUT => SYNTHESIZED_WIRE_73);


b2v_inst39 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_49,
		 Reset => SYNTHESIZED_WIRE_75,
		 dIN => SYNTHESIZED_WIRE_73,
		 ENOp => SYNTHESIZED_WIRE_52,
		 dOUT => SYNTHESIZED_WIRE_74);


b2v_inst40 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_52,
		 Reset => SYNTHESIZED_WIRE_76,
		 dIN => SYNTHESIZED_WIRE_74,
		 ENOp => SYNTHESIZED_WIRE_55,
		 dOUT => SYNTHESIZED_WIRE_75);


b2v_inst41 : delaycellv3
PORT MAP(ENp => SYNTHESIZED_WIRE_55,
		 dIN => SYNTHESIZED_WIRE_75,
		 ENOp => ENOout,
		 dOUT => SYNTHESIZED_WIRE_76);


END bdf_type;